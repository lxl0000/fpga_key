module key(
    input sys_clk,
    input sys_rst,
    input key,
    output reg key_val
);

endmodule 